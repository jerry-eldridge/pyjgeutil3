module ButterflyNet(packeti, packeto);
    input [15:0][39:0] packeti;
    output [15:0][39:0] packeto;
    reg [79:0] channel;
    reg [79:0][39:0] packetii;
    reg [79:0][39:0] packetjja;
    reg [79:0][39:0] packetjjb;
    
    assign packetii[0] = packeti[0];
    assign packetii[1] = packeti[1];
    assign packetii[2] = packeti[2];
    assign packetii[3] = packeti[3];
    assign packetii[4] = packeti[4];
    assign packetii[5] = packeti[5];
    assign packetii[6] = packeti[6];
    assign packetii[7] = packeti[7];
    assign packetii[8] = packeti[8];
    assign packetii[9] = packeti[9];
    assign packetii[10] = packeti[10];
    assign packetii[11] = packeti[11];
    assign packetii[12] = packeti[12];
    assign packetii[13] = packeti[13];
    assign packetii[14] = packeti[14];
    assign packetii[15] = packeti[15];

    ButterflyNodeD bnd000(packetii[0], channel[0]);
    ButterflyNodeD bnd001(packetii[1], channel[1]);
    ButterflyNodeD bnd002(packetii[2], channel[2]);
    ButterflyNodeD bnd003(packetii[3], channel[3]);
    ButterflyNodeD bnd004(packetii[4], channel[4]);
    ButterflyNodeD bnd005(packetii[5], channel[5]);
    ButterflyNodeD bnd006(packetii[6], channel[6]);
    ButterflyNodeD bnd007(packetii[7], channel[7]);
    ButterflyNodeD bnd008(packetii[8], channel[8]);
    ButterflyNodeD bnd009(packetii[9], channel[9]);
    ButterflyNodeD bnd010(packetii[10], channel[10]);
    ButterflyNodeD bnd011(packetii[11], channel[11]);
    ButterflyNodeD bnd012(packetii[12], channel[12]);
    ButterflyNodeD bnd013(packetii[13], channel[13]);
    ButterflyNodeD bnd014(packetii[14], channel[14]);
    ButterflyNodeD bnd015(packetii[15], channel[15]);
    ButterflyNodeD bnd016(packetii[16], channel[16]);
    ButterflyNodeD bnd017(packetii[17], channel[17]);
    ButterflyNodeD bnd018(packetii[18], channel[18]);
    ButterflyNodeD bnd019(packetii[19], channel[19]);
    ButterflyNodeD bnd020(packetii[20], channel[20]);
    ButterflyNodeD bnd021(packetii[21], channel[21]);
    ButterflyNodeD bnd022(packetii[22], channel[22]);
    ButterflyNodeD bnd023(packetii[23], channel[23]);
    ButterflyNodeD bnd024(packetii[24], channel[24]);
    ButterflyNodeD bnd025(packetii[25], channel[25]);
    ButterflyNodeD bnd026(packetii[26], channel[26]);
    ButterflyNodeD bnd027(packetii[27], channel[27]);
    ButterflyNodeD bnd028(packetii[28], channel[28]);
    ButterflyNodeD bnd029(packetii[29], channel[29]);
    ButterflyNodeD bnd030(packetii[30], channel[30]);
    ButterflyNodeD bnd031(packetii[31], channel[31]);
    ButterflyNodeD bnd032(packetii[32], channel[32]);
    ButterflyNodeD bnd033(packetii[33], channel[33]);
    ButterflyNodeD bnd034(packetii[34], channel[34]);
    ButterflyNodeD bnd035(packetii[35], channel[35]);
    ButterflyNodeD bnd036(packetii[36], channel[36]);
    ButterflyNodeD bnd037(packetii[37], channel[37]);
    ButterflyNodeD bnd038(packetii[38], channel[38]);
    ButterflyNodeD bnd039(packetii[39], channel[39]);
    ButterflyNodeD bnd040(packetii[40], channel[40]);
    ButterflyNodeD bnd041(packetii[41], channel[41]);
    ButterflyNodeD bnd042(packetii[42], channel[42]);
    ButterflyNodeD bnd043(packetii[43], channel[43]);
    ButterflyNodeD bnd044(packetii[44], channel[44]);
    ButterflyNodeD bnd045(packetii[45], channel[45]);
    ButterflyNodeD bnd046(packetii[46], channel[46]);
    ButterflyNodeD bnd047(packetii[47], channel[47]);
    ButterflyNodeD bnd048(packetii[48], channel[48]);
    ButterflyNodeD bnd049(packetii[49], channel[49]);
    ButterflyNodeD bnd050(packetii[50], channel[50]);
    ButterflyNodeD bnd051(packetii[51], channel[51]);
    ButterflyNodeD bnd052(packetii[52], channel[52]);
    ButterflyNodeD bnd053(packetii[53], channel[53]);
    ButterflyNodeD bnd054(packetii[54], channel[54]);
    ButterflyNodeD bnd055(packetii[55], channel[55]);
    ButterflyNodeD bnd056(packetii[56], channel[56]);
    ButterflyNodeD bnd057(packetii[57], channel[57]);
    ButterflyNodeD bnd058(packetii[58], channel[58]);
    ButterflyNodeD bnd059(packetii[59], channel[59]);
    ButterflyNodeD bnd060(packetii[60], channel[60]);
    ButterflyNodeD bnd061(packetii[61], channel[61]);
    ButterflyNodeD bnd062(packetii[62], channel[62]);
    ButterflyNodeD bnd063(packetii[63], channel[63]);

    switch sw000(packetii[0],channel[0], {packetjja[16],packetjjb[24]});
    switch sw001(packetii[1],channel[1], {packetjja[17],packetjjb[25]});
    switch sw002(packetii[2],channel[2], {packetjja[18],packetjjb[26]});
    switch sw003(packetii[3],channel[3], {packetjja[19],packetjjb[27]});
    switch sw004(packetii[4],channel[4], {packetjja[20],packetjjb[28]});
    switch sw005(packetii[5],channel[5], {packetjja[21],packetjjb[29]});
    switch sw006(packetii[6],channel[6], {packetjja[22],packetjjb[30]});
    switch sw007(packetii[7],channel[7], {packetjja[23],packetjjb[31]});
    switch sw008(packetii[8],channel[8], {packetjja[24],packetjjb[16]});
    switch sw009(packetii[9],channel[9], {packetjja[25],packetjjb[17]});
    switch sw010(packetii[10],channel[10], {packetjja[26],packetjjb[18]});
    switch sw011(packetii[11],channel[11], {packetjja[27],packetjjb[19]});
    switch sw012(packetii[12],channel[12], {packetjja[28],packetjjb[20]});
    switch sw013(packetii[13],channel[13], {packetjja[29],packetjjb[21]});
    switch sw014(packetii[14],channel[14], {packetjja[30],packetjjb[22]});
    switch sw015(packetii[15],channel[15], {packetjja[31],packetjjb[23]});
    switch sw016(packetii[16],channel[16], {packetjja[32],packetjjb[36]});
    switch sw017(packetii[17],channel[17], {packetjja[33],packetjjb[37]});
    switch sw018(packetii[18],channel[18], {packetjja[34],packetjjb[38]});
    switch sw019(packetii[19],channel[19], {packetjja[35],packetjjb[39]});
    switch sw020(packetii[20],channel[20], {packetjja[36],packetjjb[32]});
    switch sw021(packetii[21],channel[21], {packetjja[37],packetjjb[33]});
    switch sw022(packetii[22],channel[22], {packetjja[38],packetjjb[34]});
    switch sw023(packetii[23],channel[23], {packetjja[39],packetjjb[35]});
    switch sw024(packetii[24],channel[24], {packetjja[40],packetjjb[44]});
    switch sw025(packetii[25],channel[25], {packetjja[41],packetjjb[45]});
    switch sw026(packetii[26],channel[26], {packetjja[42],packetjjb[46]});
    switch sw027(packetii[27],channel[27], {packetjja[43],packetjjb[47]});
    switch sw028(packetii[28],channel[28], {packetjja[44],packetjjb[40]});
    switch sw029(packetii[29],channel[29], {packetjja[45],packetjjb[41]});
    switch sw030(packetii[30],channel[30], {packetjja[46],packetjjb[42]});
    switch sw031(packetii[31],channel[31], {packetjja[47],packetjjb[43]});
    switch sw032(packetii[32],channel[32], {packetjja[48],packetjjb[50]});
    switch sw033(packetii[33],channel[33], {packetjja[49],packetjjb[51]});
    switch sw034(packetii[34],channel[34], {packetjja[50],packetjjb[48]});
    switch sw035(packetii[35],channel[35], {packetjja[51],packetjjb[49]});
    switch sw036(packetii[36],channel[36], {packetjja[52],packetjjb[54]});
    switch sw037(packetii[37],channel[37], {packetjja[53],packetjjb[55]});
    switch sw038(packetii[38],channel[38], {packetjja[54],packetjjb[52]});
    switch sw039(packetii[39],channel[39], {packetjja[55],packetjjb[53]});
    switch sw040(packetii[40],channel[40], {packetjja[56],packetjjb[58]});
    switch sw041(packetii[41],channel[41], {packetjja[57],packetjjb[59]});
    switch sw042(packetii[42],channel[42], {packetjja[58],packetjjb[56]});
    switch sw043(packetii[43],channel[43], {packetjja[59],packetjjb[57]});
    switch sw044(packetii[44],channel[44], {packetjja[60],packetjjb[62]});
    switch sw045(packetii[45],channel[45], {packetjja[61],packetjjb[63]});
    switch sw046(packetii[46],channel[46], {packetjja[62],packetjjb[60]});
    switch sw047(packetii[47],channel[47], {packetjja[63],packetjjb[61]});
    switch sw048(packetii[48],channel[48], {packetjja[64],packetjjb[65]});
    switch sw049(packetii[49],channel[49], {packetjja[65],packetjjb[64]});
    switch sw050(packetii[50],channel[50], {packetjja[66],packetjjb[67]});
    switch sw051(packetii[51],channel[51], {packetjja[67],packetjjb[66]});
    switch sw052(packetii[52],channel[52], {packetjja[68],packetjjb[69]});
    switch sw053(packetii[53],channel[53], {packetjja[69],packetjjb[68]});
    switch sw054(packetii[54],channel[54], {packetjja[70],packetjjb[71]});
    switch sw055(packetii[55],channel[55], {packetjja[71],packetjjb[70]});
    switch sw056(packetii[56],channel[56], {packetjja[72],packetjjb[73]});
    switch sw057(packetii[57],channel[57], {packetjja[73],packetjjb[72]});
    switch sw058(packetii[58],channel[58], {packetjja[74],packetjjb[75]});
    switch sw059(packetii[59],channel[59], {packetjja[75],packetjjb[74]});
    switch sw060(packetii[60],channel[60], {packetjja[76],packetjjb[77]});
    switch sw061(packetii[61],channel[61], {packetjja[77],packetjjb[76]});
    switch sw062(packetii[62],channel[62], {packetjja[78],packetjjb[79]});
    switch sw063(packetii[63],channel[63], {packetjja[79],packetjjb[78]});

    assign packetii[16] = (packetjja[16]|packetjjb[16]);
    assign packetii[17] = (packetjja[17]|packetjjb[17]);
    assign packetii[18] = (packetjja[18]|packetjjb[18]);
    assign packetii[19] = (packetjja[19]|packetjjb[19]);
    assign packetii[20] = (packetjja[20]|packetjjb[20]);
    assign packetii[21] = (packetjja[21]|packetjjb[21]);
    assign packetii[22] = (packetjja[22]|packetjjb[22]);
    assign packetii[23] = (packetjja[23]|packetjjb[23]);
    assign packetii[24] = (packetjja[24]|packetjjb[24]);
    assign packetii[25] = (packetjja[25]|packetjjb[25]);
    assign packetii[26] = (packetjja[26]|packetjjb[26]);
    assign packetii[27] = (packetjja[27]|packetjjb[27]);
    assign packetii[28] = (packetjja[28]|packetjjb[28]);
    assign packetii[29] = (packetjja[29]|packetjjb[29]);
    assign packetii[30] = (packetjja[30]|packetjjb[30]);
    assign packetii[31] = (packetjja[31]|packetjjb[31]);
    assign packetii[32] = (packetjja[32]|packetjjb[32]);
    assign packetii[33] = (packetjja[33]|packetjjb[33]);
    assign packetii[34] = (packetjja[34]|packetjjb[34]);
    assign packetii[35] = (packetjja[35]|packetjjb[35]);
    assign packetii[36] = (packetjja[36]|packetjjb[36]);
    assign packetii[37] = (packetjja[37]|packetjjb[37]);
    assign packetii[38] = (packetjja[38]|packetjjb[38]);
    assign packetii[39] = (packetjja[39]|packetjjb[39]);
    assign packetii[40] = (packetjja[40]|packetjjb[40]);
    assign packetii[41] = (packetjja[41]|packetjjb[41]);
    assign packetii[42] = (packetjja[42]|packetjjb[42]);
    assign packetii[43] = (packetjja[43]|packetjjb[43]);
    assign packetii[44] = (packetjja[44]|packetjjb[44]);
    assign packetii[45] = (packetjja[45]|packetjjb[45]);
    assign packetii[46] = (packetjja[46]|packetjjb[46]);
    assign packetii[47] = (packetjja[47]|packetjjb[47]);
    assign packetii[48] = (packetjja[48]|packetjjb[48]);
    assign packetii[49] = (packetjja[49]|packetjjb[49]);
    assign packetii[50] = (packetjja[50]|packetjjb[50]);
    assign packetii[51] = (packetjja[51]|packetjjb[51]);
    assign packetii[52] = (packetjja[52]|packetjjb[52]);
    assign packetii[53] = (packetjja[53]|packetjjb[53]);
    assign packetii[54] = (packetjja[54]|packetjjb[54]);
    assign packetii[55] = (packetjja[55]|packetjjb[55]);
    assign packetii[56] = (packetjja[56]|packetjjb[56]);
    assign packetii[57] = (packetjja[57]|packetjjb[57]);
    assign packetii[58] = (packetjja[58]|packetjjb[58]);
    assign packetii[59] = (packetjja[59]|packetjjb[59]);
    assign packetii[60] = (packetjja[60]|packetjjb[60]);
    assign packetii[61] = (packetjja[61]|packetjjb[61]);
    assign packetii[62] = (packetjja[62]|packetjjb[62]);
    assign packetii[63] = (packetjja[63]|packetjjb[63]);
    assign packetii[64] = (packetjja[64]|packetjjb[64]);
    assign packetii[65] = (packetjja[65]|packetjjb[65]);
    assign packetii[66] = (packetjja[66]|packetjjb[66]);
    assign packetii[67] = (packetjja[67]|packetjjb[67]);
    assign packetii[68] = (packetjja[68]|packetjjb[68]);
    assign packetii[69] = (packetjja[69]|packetjjb[69]);
    assign packetii[70] = (packetjja[70]|packetjjb[70]);
    assign packetii[71] = (packetjja[71]|packetjjb[71]);
    assign packetii[72] = (packetjja[72]|packetjjb[72]);
    assign packetii[73] = (packetjja[73]|packetjjb[73]);
    assign packetii[74] = (packetjja[74]|packetjjb[74]);
    assign packetii[75] = (packetjja[75]|packetjjb[75]);
    assign packetii[76] = (packetjja[76]|packetjjb[76]);
    assign packetii[77] = (packetjja[77]|packetjjb[77]);
    assign packetii[78] = (packetjja[78]|packetjjb[78]);
    assign packetii[79] = (packetjja[79]|packetjjb[79]);

    assign packeto[0] = packetii[64];
    assign packeto[1] = packetii[65];
    assign packeto[2] = packetii[66];
    assign packeto[3] = packetii[67];
    assign packeto[4] = packetii[68];
    assign packeto[5] = packetii[69];
    assign packeto[6] = packetii[70];
    assign packeto[7] = packetii[71];
    assign packeto[8] = packetii[72];
    assign packeto[9] = packetii[73];
    assign packeto[10] = packetii[74];
    assign packeto[11] = packetii[75];
    assign packeto[12] = packetii[76];
    assign packeto[13] = packetii[77];
    assign packeto[14] = packetii[78];
    assign packeto[15] = packetii[79];

endmodule
